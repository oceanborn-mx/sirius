module Multiplicador_4x4 (
	input [3:0]	A,B,	//	Operandos 
	output[7:0] M		//	Producto
	);			   
	
	assign	M = A * B;
	
endmodule
