module Sumador_12b (
	input[11:0]	A,B,	//	Operandos
	output[11:0]	SUM		//	Suma
	);	 
	
	assign	SUM = A + B;
	
endmodule
